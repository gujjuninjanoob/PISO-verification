// Declaring all the required parameters
