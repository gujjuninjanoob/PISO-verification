`include "parallel_to_serial_base_test.svh"
